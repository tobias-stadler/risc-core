module CoreTB(
    input logic clk,
    input logic rst
);

endmodule
