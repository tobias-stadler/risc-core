module Top(
    input clk,
    input rst
);

endmodule
