module VivadoTop ();

  Core m_core();

endmodule
