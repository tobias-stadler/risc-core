package Mem;
  typedef logic [29:0] waddr_t;
  typedef logic [30:0] haddr_t;
  typedef logic [31:0] baddr_t;

  typedef logic [31:0] w_t;
  typedef logic [15:0] hw_t;
  typedef logic [7:0] b_t;
endpackage
